module hello;
initial 
begin
$display("hell world");
$finish;
end
endmodule